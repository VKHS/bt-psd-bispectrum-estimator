// window_fir.v
// Applies a time-domain window w[n] to incoming real samples.
// Coefficients are stored in a ROM initialized from a .mem file.
// This is a simple "one tap per sample" filter.

`ifndef WINDOW_FIR_V
`define WINDOW_FIR_V

module window_fir #(
    parameter DATA_W    = 16,
    parameter FRAC_W    = 14,
    parameter ADDR_W    = 10,              // supports up to 1024 samples
    parameter WIN_FILE  = "window_hann.mem" // generated by Python
)(
    input  wire                     clk,
    input  wire                     rst_n,
    input  wire                     in_valid,
    input  wire [ADDR_W-1:0]        in_index,   // position within frame
    input  wire signed [DATA_W-1:0] in_sample,
    output reg                      out_valid,
    output reg  signed [DATA_W-1:0] out_sample
);
    // Window coefficient ROM (Q(FRAC_W))
    reg signed [DATA_W-1:0] w_rom [0:(1<<ADDR_W)-1];

    initial begin
        $readmemh(WIN_FILE, w_rom);
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            out_valid  <= 1'b0;
            out_sample <= '0;
        end else begin
            if (in_valid) begin
                // Multiply in_sample * w[in_index] with built-in multiplier
                out_sample <= (in_sample * w_rom[in_index]) >>> FRAC_W;
                out_valid  <= 1'b1;
            end else begin
                out_valid  <= 1'b0;
            end
        end
    end
endmodule

`endif
