// cru_shared.v
// Central Rotational Unit (CRU): shared complex multiplier
// with twiddle ROM.
//
// Interface:
//  - Ready/Valid handshake on request and response.
//  - angle_idx selects twiddle e^{-j*2π*angle_idx/N_TW}.
//
// This is a "logical CRU": hardware uses a single complex multiplier
// shared between FFT, FD, window, bispectrum, etc.

`ifndef CRU_SHARED_V
`define CRU_SHARED_V

`include "complex_fixed.v"

module cru_shared #(
    parameter DATA_W   = 16,
    parameter FRAC_W   = 14,
    parameter ANGLE_W  = 9,   // e.g. 9 bits -> up to 512 twiddles
    parameter N_TW     = 512  // number of entries in twiddle ROM
)(
    input  wire                     clk,
    input  wire                     rst_n,

    // Request side
    input  wire                     req_valid,
    output wire                     req_ready,
    input  wire signed [DATA_W-1:0] xr,
    input  wire signed [DATA_W-1:0] xi,
    input  wire [ANGLE_W-1:0]       angle_idx,

    // Response side
    output reg                      resp_valid,
    input  wire                     resp_ready,
    output reg  signed [DATA_W-1:0] yr,
    output reg  signed [DATA_W-1:0] yi
);

    // Single-cycle pipeline: accept when response stage is free
    assign req_ready = (~resp_valid) | resp_ready;

    // Twiddle ROMs (cos and -sin to realize e^{-jθ})
    wire signed [DATA_W-1:0] twr;
    wire signed [DATA_W-1:0] twi;

    rom_sync #(
        .DATA_W (DATA_W),
        .ADDR_W (ANGLE_W),
        .INIT_FILE ("twiddle_cos.mem")  // generated by Python
    ) twiddle_cos_rom (
        .clk  (clk),
        .addr (angle_idx),
        .dout (twr)
    );

    rom_sync #(
        .DATA_W (DATA_W),
        .ADDR_W (ANGLE_W),
        .INIT_FILE ("twiddle_sin_neg.mem") // -sin(angle)
    ) twiddle_sin_rom (
        .clk  (clk),
        .addr (angle_idx),
        .dout (twi)
    );

    // Complex multiply using shared complex_mul block
    wire signed [DATA_W-1:0] mul_r, mul_i;

    complex_mul #(
        .DATA_W (DATA_W),
        .FRAC_W (FRAC_W)
    ) u_cmul (
        .ar (xr),
        .ai (xi),
        .br (twr),
        .bi (twi),
        .yr (mul_r),
        .yi (mul_i)
    );

    // Simple 1-stage handshake
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            resp_valid <= 1'b0;
            yr <= '0;
            yi <= '0;
        end else begin
            if (req_valid && req_ready) begin
                // Take multiply result immediately (combinational)
                yr <= mul_r;
                yi <= mul_i;
                resp_valid <= 1'b1;
            end else if (resp_valid && resp_ready) begin
                resp_valid <= 1'b0;
            end
        end
    end

endmodule


// Simple synchronous ROM for coeffs / twiddles
module rom_sync #(
    parameter DATA_W   = 16,
    parameter ADDR_W   = 9,
    parameter INIT_FILE = ""
)(
    input  wire                 clk,
    input  wire [ADDR_W-1:0]    addr,
    output reg  [DATA_W-1:0]    dout
);
    reg [DATA_W-1:0] mem [0:(1<<ADDR_W)-1];

    initial begin
        if (INIT_FILE != "") begin
            $readmemh(INIT_FILE, mem);
        end
    end

    always @(posedge clk) begin
        dout <= mem[addr];
    end
endmodule

`endif
